--   __   __     __  __     __         __
--  /\ "-.\ \   /\ \/\ \   /\ \       /\ \
--  \ \ \-.  \  \ \ \_\ \  \ \ \____  \ \ \____
--   \ \_\\"\_\  \ \_____\  \ \_____\  \ \_____\
--    \/_/ \/_/   \/_____/   \/_____/   \/_____/
--   ______     ______       __     ______     ______     ______
--  /\  __ \   /\  == \     /\ \   /\  ___\   /\  ___\   /\__  _\
--  \ \ \/\ \  \ \  __<    _\_\ \  \ \  __\   \ \ \____  \/_/\ \/
--   \ \_____\  \ \_____\ /\_____\  \ \_____\  \ \_____\    \ \_\
--    \/_____/   \/_____/ \/_____/   \/_____/   \/_____/     \/_/
--
-- https://joshbassett.info
-- https://twitter.com/nullobject
-- https://github.com/nullobject
--
-- Copyright (c) 2020 Josh Bassett
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

-- This SDRAM controller provides a symmetric 32-bit synchronous read/write
-- interface for a 16Mx16-bit SDRAM chip (e.g. AS4C16M16SA-6TCN, IS42S16400F,
-- etc.).
entity sdram is
  generic (
    -- clock frequency (in MHz)
    --
    -- This value must be provided, as it is used to calculate the number of
    -- clock cycles required for the other timing values.
    -- Both the clk and clk_in use the same frequency.
    CLK_FREQ : real;

    -- When clk_in is enabled, the clk_in signal is used for sampling the
    -- sdram_dq signal. Otherwise the clk signal is used.
    CLK_IN_ENABLE : boolean := false;

    -- 32-bit controller interface
    ADDR_WIDTH : natural := 23;
    DATA_WIDTH : natural := 32;

    -- SDRAM interface
    SDRAM_ADDR_WIDTH : natural := 13;
    SDRAM_DATA_WIDTH : natural := 16;
    SDRAM_COL_WIDTH  : natural := 9;
    SDRAM_ROW_WIDTH  : natural := 13;
    SDRAM_BANK_WIDTH : natural := 2;

    -- The delay in clock cycles, between the start of a read command and the
    -- availability of the output data.
    CAS_LATENCY : natural := 2; -- 2=below 133MHz, 3=above 133MHz

    -- The number of 16-bit words to be bursted during a read/write.
    BURST_LENGTH : natural := 2;

    -- timing values (in nanoseconds)
    --
    -- These values can be adjusted to match the exact timing of your SDRAM
    -- chip (refer to the datasheet).
    T_DESL : real := 200000.0; -- startup delay
    T_MRD  : real :=     12.0; -- mode register cycle time
    T_RC   : real :=     60.0; -- row cycle time
    T_RCD  : real :=     18.0; -- RAS to CAS delay
    T_RP   : real :=     18.0; -- precharge to activate delay
    T_WR   : real :=     12.0; -- write recovery time
    T_REFI : real :=   7800.0  -- average refresh interval
  );
  port (
    -- reset
    reset : in std_logic := '0';

    -- clock for the controller and the output signals
    clk : in std_logic;

    -- Clock for the input signals (used for sampling sdram_dq). This clock
    -- should be the same frequency as clk, but with a phase that compensates
    -- for DQ signal delay. The positive flank of this clock should coincide
    -- with the optimum DQ signal sample time.
    -- Required if CLK_IN_ENABLE is true.
    clk_in : in std_logic := 'X';

    -- address bus
    addr : in unsigned(ADDR_WIDTH-1 downto 0);

    -- input data bus
    data : in std_logic_vector(DATA_WIDTH-1 downto 0);

    -- When the write enable signal is asserted, a write operation will be performed.
    we : in std_logic;

    -- Byte select for write operations ('1' = enable byte)
    sel : in std_logic_vector(DATA_WIDTH/8-1 downto 0);

    -- When the request signal is asserted, an operation will be performed.
    req : in std_logic;

    -- The ready signal is asserted when the controller is ready to accept a
    -- new request.
    ready : out std_logic;

    -- The acknowledge signal is asserted by the SDRAM controller when
    -- a request has been accepted.
    ack : out std_logic;

    -- The valid signal is asserted when there is a valid word on the output
    -- data bus.
    valid : out std_logic;

    -- output data bus
    q : out std_logic_vector(DATA_WIDTH-1 downto 0);

    -- SDRAM interface (e.g. AS4C16M16SA-6TCN, IS42S16400F, etc.)
    sdram_a     : out unsigned(SDRAM_ADDR_WIDTH-1 downto 0);
    sdram_ba    : out unsigned(SDRAM_BANK_WIDTH-1 downto 0);
    sdram_dq    : inout std_logic_vector(SDRAM_DATA_WIDTH-1 downto 0);
    sdram_cke   : out std_logic;
    sdram_cs_n  : out std_logic;
    sdram_ras_n : out std_logic;
    sdram_cas_n : out std_logic;
    sdram_we_n  : out std_logic;
    sdram_dqm   : out std_logic_vector(SDRAM_DATA_WIDTH/8-1 downto 0)
  );
end sdram;

architecture arch of sdram is
  function ilog2(n : natural) return natural is
  begin
    return natural(ceil(log2(real(n))));
  end ilog2;

  -- Convert a ROW address to a signal suitable for sdram_a.
  function row2addr(x : unsigned) return unsigned is
  begin
    return resize(x, SDRAM_ADDR_WIDTH);
  end row2addr;

  -- Convert a COL address to a signal suitable for sdram_a.
  function col2addr(x : unsigned) return unsigned is
    variable a : unsigned(SDRAM_ADDR_WIDTH-2 downto 0);
  begin
    a := resize(x, SDRAM_ADDR_WIDTH-1);
    -- A10 = '1' -> auto precharge
    return a(SDRAM_ADDR_WIDTH-2 downto 10) & "1" & a(9 downto 0);
  end col2addr;

  -- Number of cycles that the DQ signal is delayed relative to the
  -- CAS_LATENCY cycle.
  function extra_read_latency return natural is
  begin
    if CLK_IN_ENABLE then
      -- If we use clk_in for sampling we effectively get an extra
      -- cycle of delay.
      return 1;
    else
      return 0;
    end if;
  end extra_read_latency;


  subtype command_t is std_logic_vector(3 downto 0);

  -- commands
  constant CMD_DESELECT     : command_t := "1---";
  constant CMD_LOAD_MODE    : command_t := "0000";
  constant CMD_AUTO_REFRESH : command_t := "0001";
  constant CMD_PRECHARGE    : command_t := "0010";
  constant CMD_ACTIVE       : command_t := "0011";
  constant CMD_WRITE        : command_t := "0100";
  constant CMD_READ         : command_t := "0101";
  constant CMD_STOP         : command_t := "0110";
  constant CMD_NOP          : command_t := "0111";

  -- the ordering of the accesses within a burst
  constant BURST_TYPE : std_logic := '0'; -- 0=sequential, 1=interleaved

  -- the write burst mode enables bursting for write operations
  constant WRITE_BURST_MODE : std_logic := '0'; -- 0=burst, 1=single

  -- the value written to the address bus during initialization
  constant INIT_CMD : unsigned(SDRAM_ADDR_WIDTH-1 downto 0) := (
    to_unsigned(0, SDRAM_ADDR_WIDTH-11) &
    "10000000000"
  );

  -- the value written to the mode register to configure the memory
  constant MODE_REG : unsigned(SDRAM_ADDR_WIDTH-1 downto 0) := (
    to_unsigned(0, SDRAM_ADDR_WIDTH-10) &
    WRITE_BURST_MODE &
    "00" &
    to_unsigned(CAS_LATENCY, 3) &
    BURST_TYPE &
    to_unsigned(ilog2(BURST_LENGTH), 3)
  );

  -- calculate the clock period (in nanoseconds)
  constant CLK_PERIOD : real := 1.0/CLK_FREQ*1000.0;

  -- the number of clock cycles to wait before initialising the device
  constant INIT_WAIT : natural := natural(ceil(T_DESL/CLK_PERIOD));

  -- the number of clock cycles to wait while a LOAD MODE command is being
  -- executed
  constant LOAD_MODE_WAIT : natural := natural(ceil(T_MRD/CLK_PERIOD));

  -- the number of clock cycles to wait while an ACTIVE command is being
  -- executed
  constant ACTIVE_WAIT : natural := natural(ceil(T_RCD/CLK_PERIOD));

  -- the number of clock cycles to wait while a REFRESH command is being
  -- executed
  constant REFRESH_WAIT : natural := natural(ceil(T_RC/CLK_PERIOD));

  -- the number of clock cycles to wait while a PRECHARGE command is being
  -- executed
  constant PRECHARGE_WAIT : natural := natural(ceil(T_RP/CLK_PERIOD));

  -- the number of clock cycles to wait while a READ command is being executed
  constant READ_WAIT : natural := CAS_LATENCY+BURST_LENGTH;

  -- the number of clock cycles to wait while a WRITE command is being executed
  constant WRITE_WAIT : natural := BURST_LENGTH+natural(ceil((T_WR+T_RP)/CLK_PERIOD));

  -- the number of clock cycles before the memory controller needs to refresh
  -- the SDRAM
  constant REFRESH_INTERVAL : natural := natural(floor(T_REFI/CLK_PERIOD))-10;

  type state_t is (INIT, MODE, IDLE, ACTIVE, READ, WRITE, REFRESH);

  -- state signals
  signal state, next_state : state_t;

  -- command signals
  signal cmd, next_cmd : command_t := CMD_NOP;

  -- control signals
  signal start          : std_logic;
  signal load_mode_done : std_logic;
  signal active_done    : std_logic;
  signal refresh_done   : std_logic;
  signal read_done      : std_logic;
  signal write_done     : std_logic;
  signal should_refresh : std_logic;

  -- counters
  constant MAX_WAIT_COUNT    : natural := INIT_WAIT+PRECHARGE_WAIT+REFRESH_WAIT+REFRESH_WAIT+1;
  constant MAX_REFRESH_COUNT : natural := REFRESH_INTERVAL;
  signal wait_counter    : natural range 0 to MAX_WAIT_COUNT;
  signal refresh_counter : natural range 0 to MAX_REFRESH_COUNT;

  -- registers
  signal addr_reg  : unsigned(SDRAM_COL_WIDTH+SDRAM_ROW_WIDTH+SDRAM_BANK_WIDTH-1 downto 0);
  signal data_reg  : std_logic_vector(DATA_WIDTH-1 downto 0);
  signal we_reg    : std_logic;
  signal sel_n_reg : std_logic_vector(DATA_WIDTH/8-1 downto 0);
  signal q_reg     : std_logic_vector(DATA_WIDTH-1 downto 0);

  -- DQ signal, sampled in the clk_in clock domain
  signal dq_in : std_logic_vector(SDRAM_DATA_WIDTH-1 downto 0);

  -- aliases to decode the address register
  alias col  : unsigned(SDRAM_COL_WIDTH-1 downto 0) is addr_reg(SDRAM_COL_WIDTH-1 downto 0);
  alias row  : unsigned(SDRAM_ROW_WIDTH-1 downto 0) is addr_reg(SDRAM_COL_WIDTH+SDRAM_ROW_WIDTH-1 downto SDRAM_COL_WIDTH);
  alias bank : unsigned(SDRAM_BANK_WIDTH-1 downto 0) is addr_reg(SDRAM_COL_WIDTH+SDRAM_ROW_WIDTH+SDRAM_BANK_WIDTH-1 downto SDRAM_COL_WIDTH+SDRAM_ROW_WIDTH);
begin
  -- state machine
  fsm : process (state, wait_counter, req, we_reg, sel_n_reg, load_mode_done, active_done, refresh_done, read_done, write_done, should_refresh)
  begin
    next_state <= state;

    -- default to a NOP command
    next_cmd <= CMD_NOP;

    case state is
      -- execute the initialisation sequence
      when INIT =>
        if wait_counter = 0 then
          next_cmd <= CMD_DESELECT;
        elsif wait_counter = INIT_WAIT-1 then
          next_cmd <= CMD_PRECHARGE;
        elsif wait_counter = INIT_WAIT+PRECHARGE_WAIT-1 then
          next_cmd <= CMD_AUTO_REFRESH;
        elsif wait_counter = INIT_WAIT+PRECHARGE_WAIT+REFRESH_WAIT-1 then
          next_cmd <= CMD_AUTO_REFRESH;
        elsif wait_counter = INIT_WAIT+PRECHARGE_WAIT+REFRESH_WAIT+REFRESH_WAIT-1 then
          next_state <= MODE;
          next_cmd   <= CMD_LOAD_MODE;
        end if;

      -- load the mode register
      when MODE =>
        if load_mode_done = '1' then
          next_state <= IDLE;
        end if;

      -- wait for a read/write request
      when IDLE =>
        if should_refresh = '1' then
          next_state <= REFRESH;
          next_cmd   <= CMD_AUTO_REFRESH;
        elsif req = '1' then
          next_state <= ACTIVE;
          next_cmd   <= CMD_ACTIVE;
        end if;

      -- activate the row
      when ACTIVE =>
        if active_done = '1' then
          if we_reg = '1' then
            next_state <= WRITE;
            next_cmd   <= CMD_WRITE;
          else
            next_state <= READ;
            next_cmd   <= CMD_READ;
          end if;
        end if;

      -- execute a read command
      when READ =>
        if read_done = '1' then
          if should_refresh = '1' then
            next_state <= REFRESH;
            next_cmd   <= CMD_AUTO_REFRESH;
          elsif req = '1' then
            next_state <= ACTIVE;
            next_cmd   <= CMD_ACTIVE;
          else
            next_state <= IDLE;
          end if;
        end if;

      -- execute a write command
      when WRITE =>
        if write_done = '1' then
          if should_refresh = '1' then
            next_state <= REFRESH;
            next_cmd   <= CMD_AUTO_REFRESH;
          elsif req = '1' then
            next_state <= ACTIVE;
            next_cmd   <= CMD_ACTIVE;
          else
            next_state <= IDLE;
          end if;
        end if;

      -- execute an auto refresh
      when REFRESH =>
        if refresh_done = '1' then
          if req = '1' then
            next_state <= ACTIVE;
            next_cmd   <= CMD_ACTIVE;
          else
            next_state <= IDLE;
          end if;
        end if;
    end case;
  end process;

  -- latch the next state
  latch_next_state : process (clk, reset)
  begin
    if reset = '1' then
      state <= INIT;
      cmd   <= CMD_NOP;
    elsif rising_edge(clk) then
      state <= next_state;
      cmd   <= next_cmd;
    end if;
  end process;

  -- the wait counter is used to hold the current state for a number of clock
  -- cycles
  update_wait_counter : process (clk, reset)
  begin
    if reset = '1' then
      wait_counter <= 0;
    elsif rising_edge(clk) then
      if state /= next_state then -- state changing
        wait_counter <= 0;
      elsif state = IDLE then    -- counter would overflow when IDLE
        wait_counter <= 0;
      else
        wait_counter <= wait_counter + 1;
      end if;
    end if;
  end process;

  -- the refresh counter is used to periodically trigger a refresh operation
  update_refresh_counter : process (clk, reset)
  begin
    if reset = '1' then
      refresh_counter <= 0;
    elsif rising_edge(clk) then
      if state = REFRESH and wait_counter = 0 then
        refresh_counter <= 0;
      elsif refresh_counter /= MAX_REFRESH_COUNT then
        refresh_counter <= refresh_counter + 1;
      end if;
    end if;
  end process;

  -- latch the rquest
  latch_request : process (reset, clk)
  begin
    if reset = '1' then
      addr_reg <= (others => '0');
      data_reg <= (others => '0');
      we_reg <= '0';
      sel_n_reg <= (others => '0');
    elsif rising_edge(clk) then
      if start = '1' then
        -- we need to multiply the address by two, because we are converting
        -- from a 32-bit controller address to a 16-bit SDRAM address
        addr_reg  <= shift_left(resize(addr, addr_reg'length), 1);
        data_reg  <= data;
        we_reg    <= we;
        sel_n_reg <= not sel;
      end if;
    end if;
  end process;

  -- set wait signals
  load_mode_done <= '1' when wait_counter = LOAD_MODE_WAIT-1 else '0';
  active_done    <= '1' when wait_counter = ACTIVE_WAIT-1    else '0';
  refresh_done   <= '1' when wait_counter = REFRESH_WAIT-1   else '0';
  read_done      <= '1' when wait_counter = READ_WAIT-1      else '0';
  write_done     <= '1' when wait_counter = WRITE_WAIT-1     else '0';

  -- the SDRAM should be refreshed when the refresh interval has elapsed
  should_refresh <= '1' when refresh_counter >= REFRESH_INTERVAL-1 else '0';

  -- a new request is only allowed at the end of the IDLE, READ, WRITE, and
  -- REFRESH states
  start <= '1' when (state = IDLE) or
                    (state = READ and read_done = '1') or
                    (state = WRITE and write_done = '1') or
                    (state = REFRESH and refresh_done = '1') else '0';

  -- assert the ready signal when we're ready to accept a new request
  ready <= start;

  -- assert the acknowledge signal at the beginning of the ACTIVE state
  ack <= '1' when state = ACTIVE and wait_counter = 0 else '0';

  -- set output data
  q <= q_reg;

  -- deassert the clock enable at the beginning of the INIT state
  sdram_cke <= '0' when state = INIT and wait_counter = 0 else '1';

  -- set SDRAM control signals
  (sdram_cs_n, sdram_ras_n, sdram_cas_n, sdram_we_n) <= cmd;

  -- set SDRAM bank
  with state select
    sdram_ba <=
      bank            when ACTIVE,
      bank            when READ,
      bank            when WRITE,
      (others => '0') when others;

  -- set SDRAM address
  with state select
    sdram_a <=
      INIT_CMD        when INIT,
      MODE_REG        when MODE,
      row2addr(row)   when ACTIVE,
      col2addr(col)   when READ,
      col2addr(col)   when WRITE,
      (others => '0') when others;

  DQ_IN_GEN : if CLK_IN_ENABLE generate
    -- This is a FF that latches the DQ signal in the clk_in clock domain.
    process (reset, clk_in)
    begin
      if reset = '1' then
        dq_in <= (others => '0');
      elsif rising_edge(clk_in) then
        dq_in <= sdram_dq;
      end if;
    end process;
  else generate
    -- Just forward the sdram_dq signal without a FF.
    dq_in <= sdram_dq;
  end generate;

  -- read the next sub-word as it's bursted from the SDRAM
  process (reset, clk)
    constant C_MAX_BURST_CNT : natural := BURST_LENGTH + extra_read_latency;
    variable v_burst_cnt : natural range 0 to C_MAX_BURST_CNT := C_MAX_BURST_CNT;
    variable v_idx : natural;
  begin
    if reset = '1' then
      q_reg <= (others => '0');
      valid <= '0';
    elsif rising_edge(clk) then
      -- Which sub-word are we currently reading?
      if state = READ and wait_counter = CAS_LATENCY then
        v_burst_cnt := 0;
      elsif v_burst_cnt < C_MAX_BURST_CNT then
        v_burst_cnt := v_burst_cnt + 1;
      end if;

      if v_burst_cnt >= extra_read_latency and v_burst_cnt < C_MAX_BURST_CNT then
        v_idx := v_burst_cnt - extra_read_latency;
        q_reg(SDRAM_DATA_WIDTH*(v_idx+1)-1 downto SDRAM_DATA_WIDTH*v_idx) <= dq_in;
      end if;

      -- Was this the final sub-word?
      if v_burst_cnt = (C_MAX_BURST_CNT - 1) then
        valid <= '1';
      else
        valid <= '0';
      end if;
    end if;
  end process;

  -- write the next sub-word from the write buffer
  process (data_reg, sel_n_reg, state, wait_counter)
  begin
    -- TODO(m): Add support for other DATA_WIDTH/BURST_LENGTH/etc settings.
    if state = WRITE and wait_counter = 0 then
      sdram_dq <= data_reg(SDRAM_DATA_WIDTH-1 downto 0);
      sdram_dqm(1) <= sel_n_reg(1);
      sdram_dqm(0) <= sel_n_reg(0);
    elsif state = WRITE and wait_counter = 1 then
      sdram_dq <= data_reg(SDRAM_DATA_WIDTH*2-1 downto SDRAM_DATA_WIDTH);
      sdram_dqm(1) <= sel_n_reg(3);
      sdram_dqm(0) <= sel_n_reg(2);
    else
      sdram_dq <= (others => 'Z');
      sdram_dqm(1) <= '0';
      sdram_dqm(0) <= '0';
    end if;
  end process;
end architecture arch;
